// Code your design here
module or_(a,b,c);
  input a,b;
  output c;
  assign c=a | b;
endmodule